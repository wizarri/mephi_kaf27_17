module tausworthe_mod
(
  input clk, rst,clk_lr,
  output [31:0] generator_out
);
  wire [31:0] out1, out2, out3;
  tausworthe
  #(
  	.SEED(32'hE761B9DB), .CONST(32'hE4B4D358), 
  	.SHIFT_L1(8'd13), .SHIFT_L2(8'd12), .SHIFT_R(8'd19)
  )
  part_1
  (
    .clk(clk),
	 .clk_lr(clk_lr),
    .rst(rst),
    .out(out1) 
  );

  tausworthe 
  #(
  	.SEED(32'hB4B4D15C), .CONST(32'h84B4D155), 
  	.SHIFT_L1(4'd2), .SHIFT_L2(4'd4), .SHIFT_R(8'd25)
  )
  part_2
  (
    .clk(clk),
	 .clk_lr(clk_lr),
    .rst(rst),
    .out(out2) 
  );

  tausworthe 
  #(
  	.SEED(32'hC0B4DD55), .CONST(32'h86B4C155), 
  	.SHIFT_L1(4'd3), .SHIFT_L2(8'd17), .SHIFT_R(8'd11)
  )
  part_3
  (
    .clk(clk),
	 .clk_lr(clk_lr),
    .rst(rst),
    .out(out3) 
  );

  assign generator_out = out1 ^ out2 ^ out3;

endmodule // tausworthe