модуль  hello_world ();
input i0 // YRR
input i1 // YRR
endmodule